`ifndef __DEFINE_V
`define __DEFINE_V

`include "config.sv"

`define AVALON_BURST_COUNT_WIDTH          (8)

`endif