module core_ma_lsu (
  ports
);
  
endmodule