`ifndef __CONFIG_V
`define __CONFIG_V

/****************************************************************************************
选择FPGA类型,将通过该选项对内部的RAM进行适配
可选项：
	FPGA_TYPE_ALTERA
	FPGA_TYPE_XILINX
	FPGA_TYPE_NULL
****************************************************************************************/
`define FPGA_TYPE_ALTERA


/****************************************************************************************
选择FPGA复位电平
可选项：
	FPGA_REST_LEVEL_H
	FPGA_REST_LEVEL_L
****************************************************************************************/
`define FPGA_REST_LEVEL_H

`endif
