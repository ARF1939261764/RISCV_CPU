module istr_c2i (
  input[15:0]  istr_c,
  output[31:0] istr_i
);

assign istr_i=32'hFFFFFFFF;

endmodule
