module istr_c2i (
  input[15:0]  istr_c,
  output[31:0] istr_i
);



endmodule
