`ifndef __DEFINE_V
`define __DEFINE_V

`include "../config/config.sv"

`define AVALON_BURST_COUNT_WIDTH          (8)

`endif