module core();

endmodule
