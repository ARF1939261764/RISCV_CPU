module core(
  input logic clk,
  input logic rest
  
);

endmodule
