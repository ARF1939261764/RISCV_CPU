module core_if(
  input clk,
  input rest,
  
);



endmodule
