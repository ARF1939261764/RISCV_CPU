module core_ex_alu_mul_div(
  input  logic       clk,
  input  logic       rest,
  input  logic       sig,  
  input  logic[31:0] in1,
  input  logic[31:0] in2,
  output logic[63:0] out
);
  
endmodule