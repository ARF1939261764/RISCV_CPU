module avl_bus_ns2m_controller(

);

endmodule
